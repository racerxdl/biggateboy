module top (
  input  wire clk
  output memAddress[15:0],
  inout  memData[7:0]
);

// CPU Registers
reg [15:0] regPC; // Program Counter
reg [15:0] regSP; // Stack Pointer

reg [7:0] regA;
reg [7:0] regB;
reg [7:0] regC;
reg [7:0] regD;
reg [7:0] regE;

reg [7:0] regF; // Flag Register
reg [7:0] regH;
reg [7:0] regL;

wire regHL = {regH, regL};
wire regBC = {regB, regC};
wire regDE = {regD, regE};
wire regZ  = regF[7];
wire regS  = regF[6];
wire regH  = regF[5];
wire regC  = regF[4];

endmodule